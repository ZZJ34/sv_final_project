import uvm_pkg::*; 

`include "uvm_macros.svh"

`include "./interface/apb_uart_interface.sv"

`include "./object/transaction.sv"

`include "./object/sequence/base_sequence.sv"

`include "./reg_model/reg_model.sv"

`include "./component/apb_input_driver.sv"
`include "./component/apb_input_monitor.sv"
`include "./component/uart_output_monitor.sv"
`include "./component/sequencer.sv"
`include "./component/input_agent.sv"
`include "./component/output_agent.sv"
`include "./component/model.sv"
`include "./component/scoreboard.sv"
`include "./component/environment.sv"