import uvm_pkg::*; 

`include "uvm_macros.svh"

`include "./interface/apb_uart_interface.sv"

`include "./object/apb_transaction.sv"
`include "./object/uart_transaction.sv"

`include "./component/apb_input_driver.sv"
`include "./component/apb_input_monitor.sv"
`include "./component/environment.sv"